magic
tech sky130A
magscale 1 2
timestamp 1757899848
<< checkpaint >>
rect -3722 40702 35502 48552
rect -3722 -2912 67812 40702
rect 28588 -10762 67812 -2912
<< error_s >>
rect 2660 15870 2760 15945
rect 2670 15810 2820 15865
rect 20444 15178 20502 15378
rect 19198 14834 19712 14892
rect 19972 14834 20372 14892
rect 19198 14376 19712 14434
rect 19972 14376 20372 14434
rect 19198 14154 19712 14212
rect 19972 14154 20372 14212
rect 19198 13696 19712 13754
rect 19972 13696 20372 13754
rect 19198 13468 19712 13526
rect 19972 13454 20372 13512
rect 19198 13010 19712 13068
rect 19972 12996 20372 13054
rect 19198 12782 19712 12840
rect 19972 12774 20372 12832
rect 17755 12324 18450 12382
rect 18712 12324 19712 12382
rect 19972 12316 20372 12374
rect 17755 12096 18450 12154
rect 18712 12096 19712 12154
rect 19972 12094 20372 12152
rect 17755 11638 18450 11696
rect 18712 11638 19712 11696
rect 19972 11636 20372 11694
rect 17755 11414 18452 11472
rect 18712 11414 19712 11472
rect 19972 11414 20372 11472
rect 17755 10956 18452 11014
rect 18712 10956 19712 11014
rect 19972 10956 20372 11014
rect 13488 9827 13888 9885
rect 14143 9829 15143 9887
rect 15377 9830 16377 9888
rect 16630 9830 17167 9888
rect 13488 9369 13888 9427
rect 14143 9371 15143 9429
rect 15377 9372 16377 9430
rect 13488 9145 13888 9203
rect 14141 9145 15141 9203
rect 15382 9144 16382 9202
rect 13488 8687 13888 8745
rect 14141 8687 15141 8745
rect 15382 8686 16382 8744
rect 13489 8464 13889 8522
rect 14142 8464 15142 8522
rect 15381 8465 16381 8523
rect 13489 8006 13889 8064
rect 14142 8006 15142 8064
rect 15381 8007 16381 8065
<< nwell >>
rect 20530 15370 20590 15460
<< pwell >>
rect 13330 9830 13420 9920
rect 13310 5850 13440 5940
<< psubdiff >>
rect 13340 9950 13380 9974
rect 13340 9866 13380 9890
rect 13320 5920 13360 5944
rect 13320 5826 13360 5850
<< nsubdiff >>
rect 20530 15390 20550 15460
rect 20530 15370 20590 15390
<< psubdiffcont >>
rect 13340 9890 13380 9950
rect 13320 5850 13360 5920
<< nsubdiffcont >>
rect 20550 15390 20590 15460
<< locali >>
rect 20530 15390 20550 15460
rect 20530 15370 20590 15390
rect 13340 9950 13380 9966
rect 13340 9874 13380 9890
rect 13320 5920 13360 5936
rect 13320 5834 13360 5850
<< viali >>
rect 20550 15390 20590 15460
rect 13340 9890 13380 9950
rect 13320 5850 13360 5920
<< metal1 >>
rect 20530 15420 20550 15460
rect 20490 15390 20550 15420
rect 20590 15390 20600 15420
rect 20490 15340 20600 15390
rect 13330 9950 13420 9960
rect 13330 9890 13340 9950
rect 13380 9890 13420 9950
rect 13330 9830 13420 9890
rect 13310 5920 13440 6010
rect 13310 5850 13320 5920
rect 13360 5850 13440 5920
rect 13310 5840 13370 5850
<< metal3 >>
rect 27220 45022 27310 45040
rect 27220 44958 27233 45022
rect 27297 44958 27310 45022
rect 27220 44940 27310 44958
rect 27760 44950 27850 44960
rect 27760 44947 31565 44950
rect 7890 44847 8560 44870
rect 7890 44783 7948 44847
rect 8012 44783 8148 44847
rect 8212 44783 8338 44847
rect 8402 44783 8560 44847
rect 7890 44190 8560 44783
rect 27220 44800 27300 44940
rect 27760 44883 27773 44947
rect 27837 44937 31565 44947
rect 27837 44883 31478 44937
rect 27760 44873 31478 44883
rect 31542 44880 31565 44937
rect 31542 44873 31570 44880
rect 27760 44870 31570 44873
rect 31450 44827 31570 44870
rect 31130 44800 31390 44810
rect 27220 44797 31390 44800
rect 27220 44733 31158 44797
rect 31222 44787 31390 44797
rect 31222 44733 31298 44787
rect 27220 44723 31298 44733
rect 31362 44723 31390 44787
rect 31450 44763 31478 44827
rect 31542 44763 31570 44827
rect 31450 44750 31570 44763
rect 27220 44720 31390 44723
rect 31270 44710 31390 44720
rect 800 36207 2150 36220
rect 800 36143 833 36207
rect 897 36143 973 36207
rect 1037 36143 1113 36207
rect 1177 36143 2150 36207
rect 800 36087 2150 36143
rect 800 36023 833 36087
rect 897 36023 973 36087
rect 1037 36023 1113 36087
rect 1177 36023 2150 36087
rect 800 36010 2150 36023
rect 200 20977 2150 20990
rect 200 20913 233 20977
rect 297 20913 353 20977
rect 417 20913 483 20977
rect 547 20913 2150 20977
rect 200 20867 2150 20913
rect 200 20803 213 20867
rect 277 20803 343 20867
rect 407 20803 473 20867
rect 537 20803 2150 20867
rect 200 20790 2150 20803
rect 2660 15780 2760 15910
rect 21570 4937 30950 4950
rect 21570 4873 21598 4937
rect 21662 4873 21678 4937
rect 21742 4873 30778 4937
rect 30842 4873 30858 4937
rect 30922 4873 30950 4937
rect 21570 4827 30950 4873
rect 21570 4763 21598 4827
rect 21662 4763 21678 4827
rect 21742 4763 30778 4827
rect 30842 4763 30858 4827
rect 30922 4763 30950 4827
rect 21570 4750 30950 4763
rect 14906 3192 15086 3210
rect 14906 3128 14923 3192
rect 14987 3128 15003 3192
rect 15067 3128 15086 3192
rect 14906 2637 15086 3128
rect 14906 2573 14923 2637
rect 14987 2573 15003 2637
rect 15067 2573 15086 2637
rect 14906 2537 15086 2573
rect 14906 2473 14923 2537
rect 14987 2473 15003 2537
rect 15067 2473 15086 2537
rect 14906 2459 15086 2473
rect 220 1467 290 1470
rect 220 1403 223 1467
rect 287 1403 290 1467
rect 220 1400 290 1403
rect 350 1467 420 1470
rect 350 1403 353 1467
rect 417 1403 420 1467
rect 350 1400 420 1403
rect 480 1467 550 1470
rect 480 1403 483 1467
rect 547 1403 550 1467
rect 480 1400 550 1403
rect 220 1357 290 1360
rect 220 1293 223 1357
rect 287 1293 290 1357
rect 220 1290 290 1293
rect 350 1357 420 1360
rect 350 1293 353 1357
rect 417 1293 420 1357
rect 350 1290 420 1293
rect 480 1357 550 1360
rect 480 1293 483 1357
rect 547 1293 550 1357
rect 480 1290 550 1293
rect 800 1177 1200 1190
rect 800 1113 823 1177
rect 887 1113 963 1177
rect 1027 1113 1093 1177
rect 1157 1113 1200 1177
rect 800 1077 1200 1113
rect 800 1013 823 1077
rect 887 1013 963 1077
rect 1027 1013 1093 1077
rect 1157 1013 1200 1077
rect 800 1000 1200 1013
rect 800 987 21770 1000
rect 800 923 21598 987
rect 21662 923 21678 987
rect 21742 923 21770 987
rect 800 877 21770 923
rect 800 813 21598 877
rect 21662 813 21678 877
rect 21742 813 21770 877
rect 800 800 21770 813
<< via3 >>
rect 27233 44958 27297 45022
rect 7948 44783 8012 44847
rect 8148 44783 8212 44847
rect 8338 44783 8402 44847
rect 27773 44883 27837 44947
rect 31478 44873 31542 44937
rect 31158 44733 31222 44797
rect 31298 44723 31362 44787
rect 31478 44763 31542 44827
rect 833 36143 897 36207
rect 973 36143 1037 36207
rect 1113 36143 1177 36207
rect 833 36023 897 36087
rect 973 36023 1037 36087
rect 1113 36023 1177 36087
rect 233 20913 297 20977
rect 353 20913 417 20977
rect 483 20913 547 20977
rect 213 20803 277 20867
rect 343 20803 407 20867
rect 473 20803 537 20867
rect 21598 4873 21662 4937
rect 21678 4873 21742 4937
rect 30778 4873 30842 4937
rect 30858 4873 30922 4937
rect 21598 4763 21662 4827
rect 21678 4763 21742 4827
rect 30778 4763 30842 4827
rect 30858 4763 30922 4827
rect 14923 3128 14987 3192
rect 15003 3128 15067 3192
rect 14923 2573 14987 2637
rect 15003 2573 15067 2637
rect 14923 2473 14987 2537
rect 15003 2473 15067 2537
rect 223 1403 287 1467
rect 353 1403 417 1467
rect 483 1403 547 1467
rect 223 1293 287 1357
rect 353 1293 417 1357
rect 483 1293 547 1357
rect 823 1113 887 1177
rect 963 1113 1027 1177
rect 1093 1113 1157 1177
rect 823 1013 887 1077
rect 963 1013 1027 1077
rect 1093 1013 1157 1077
rect 21598 923 21662 987
rect 21678 923 21742 987
rect 21598 813 21662 877
rect 21678 813 21742 877
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 45040 27170 45152
rect 27662 45040 27722 45152
rect 27110 45022 27310 45040
rect 27110 44958 27233 45022
rect 27297 44958 27310 45022
rect 27110 44952 27310 44958
rect 27662 44960 27840 45040
rect 27662 44952 27850 44960
rect 800 44847 26647 44952
rect 27220 44940 27310 44952
rect 27760 44947 27850 44952
rect 27760 44883 27773 44947
rect 27837 44883 27850 44947
rect 28214 44938 28274 45152
rect 28766 44938 28826 45152
rect 29318 44952 29378 45152
rect 29310 44938 29378 44952
rect 27760 44870 27850 44883
rect 28210 44870 29378 44938
rect 31450 44937 31570 44950
rect 31450 44873 31478 44937
rect 31542 44873 31570 44937
rect 800 44783 7948 44847
rect 8012 44783 8148 44847
rect 8212 44783 8338 44847
rect 8402 44783 26647 44847
rect 800 44760 26647 44783
rect 28210 44760 28290 44870
rect 31450 44827 31570 44873
rect 200 20977 600 44152
rect 200 20913 233 20977
rect 297 20913 353 20977
rect 417 20913 483 20977
rect 547 20913 600 20977
rect 200 20867 600 20913
rect 200 20803 213 20867
rect 277 20803 343 20867
rect 407 20803 473 20867
rect 537 20803 600 20867
rect 200 1467 600 20803
rect 200 1403 223 1467
rect 287 1403 353 1467
rect 417 1403 483 1467
rect 547 1403 600 1467
rect 200 1357 600 1403
rect 200 1293 223 1357
rect 287 1293 353 1357
rect 417 1293 483 1357
rect 547 1293 600 1357
rect 200 1000 600 1293
rect 800 36207 1200 44760
rect 26550 44680 28290 44760
rect 31130 44797 31390 44810
rect 31130 44733 31158 44797
rect 31222 44787 31390 44797
rect 31222 44733 31298 44787
rect 31130 44723 31298 44733
rect 31362 44723 31390 44787
rect 31130 44720 31390 44723
rect 800 36143 833 36207
rect 897 36143 973 36207
rect 1037 36143 1113 36207
rect 1177 36143 1200 36207
rect 800 36087 1200 36143
rect 800 36023 833 36087
rect 897 36023 973 36087
rect 1037 36023 1113 36087
rect 1177 36023 1200 36087
rect 800 1177 1200 36023
rect 31270 15930 31390 44720
rect 31450 44763 31478 44827
rect 31542 44763 31570 44827
rect 31450 15910 31570 44763
rect 20550 15390 20590 15460
rect 22470 5210 22650 5520
rect 21100 5030 22650 5210
rect 14920 3192 15070 3200
rect 14920 3128 14923 3192
rect 14987 3128 15003 3192
rect 15067 3128 15070 3192
rect 14920 3120 15070 3128
rect 800 1113 823 1177
rect 887 1113 963 1177
rect 1027 1113 1093 1177
rect 1157 1113 1200 1177
rect 800 1077 1200 1113
rect 800 1013 823 1077
rect 887 1013 963 1077
rect 1027 1013 1093 1077
rect 1157 1013 1200 1077
rect 800 1000 1200 1013
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 2990
rect 14906 2637 15086 2650
rect 14906 2573 14923 2637
rect 14987 2573 15003 2637
rect 15067 2573 15086 2637
rect 14906 2537 15086 2573
rect 14906 2473 14923 2537
rect 14987 2473 15003 2537
rect 15067 2473 15086 2537
rect 14906 0 15086 2473
rect 21100 1540 21280 5030
rect 18770 1360 21280 1540
rect 21570 4937 21770 4950
rect 21570 4873 21598 4937
rect 21662 4873 21678 4937
rect 21742 4873 21770 4937
rect 21570 4827 21770 4873
rect 21570 4763 21598 4827
rect 21662 4763 21678 4827
rect 21742 4763 21770 4827
rect 18770 0 18950 1360
rect 21570 987 21770 4763
rect 23750 4500 23930 5670
rect 21570 923 21598 987
rect 21662 923 21678 987
rect 21742 923 21770 987
rect 21570 877 21770 923
rect 21570 813 21598 877
rect 21662 813 21678 877
rect 21742 813 21770 877
rect 21570 800 21770 813
rect 22634 4320 23930 4500
rect 24360 4560 24540 5640
rect 30750 4937 30950 4950
rect 30750 4873 30778 4937
rect 30842 4873 30858 4937
rect 30922 4873 30950 4937
rect 30750 4827 30950 4873
rect 30750 4763 30778 4827
rect 30842 4763 30858 4827
rect 30922 4763 30950 4827
rect 30750 4750 30950 4763
rect 31020 4620 31200 4970
rect 24360 4380 26678 4560
rect 22634 0 22814 4320
rect 26498 0 26678 4380
rect 30362 4440 31200 4620
rect 30362 0 30542 4440
use Diff_Opamp  Diff_Opamp_0
timestamp 1757899188
transform 0 -1 31380 1 0 4920
box -3900 -190 39700 31170
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 600 44152 1 FreeSans 500 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 500 0 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
