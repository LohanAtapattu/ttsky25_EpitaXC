magic
tech sky130A
magscale 1 2
timestamp 1757892507
<< metal3 >>
rect 27220 45030 27310 45040
rect 27220 44950 27230 45030
rect 27300 44950 27310 45030
rect 27220 44940 27310 44950
rect 27760 44950 27850 44960
rect 7890 44860 8560 44870
rect 7890 44770 7920 44860
rect 8040 44770 8120 44860
rect 8240 44770 8310 44860
rect 8430 44770 8560 44860
rect 7890 44190 8560 44770
rect 27220 44800 27300 44940
rect 27760 44880 27770 44950
rect 27840 44940 31565 44950
rect 27840 44880 31460 44940
rect 27760 44870 31460 44880
rect 31560 44880 31565 44940
rect 31560 44870 31570 44880
rect 31450 44830 31570 44870
rect 31130 44800 31390 44810
rect 27220 44730 31140 44800
rect 31240 44790 31390 44800
rect 31240 44730 31280 44790
rect 27220 44720 31280 44730
rect 31380 44720 31390 44790
rect 31450 44760 31460 44830
rect 31560 44760 31570 44830
rect 31450 44750 31570 44760
rect 31270 44710 31390 44720
rect 800 36210 2150 36220
rect 800 36140 820 36210
rect 910 36140 960 36210
rect 1050 36140 1100 36210
rect 1190 36140 2150 36210
rect 800 36090 2150 36140
rect 800 36020 820 36090
rect 910 36020 960 36090
rect 1050 36020 1100 36090
rect 1190 36020 2150 36090
rect 800 36010 2150 36020
rect 200 20980 2150 20990
rect 200 20910 230 20980
rect 300 20910 350 20980
rect 420 20910 480 20980
rect 550 20910 2150 20980
rect 200 20870 2150 20910
rect 200 20800 210 20870
rect 280 20800 340 20870
rect 410 20800 470 20870
rect 540 20800 2150 20870
rect 200 20790 2150 20800
rect 21570 4940 30950 4950
rect 21570 4870 21590 4940
rect 21750 4870 30760 4940
rect 30940 4870 30950 4940
rect 21570 4830 30950 4870
rect 21570 4760 21590 4830
rect 21750 4760 30760 4830
rect 30940 4760 30950 4830
rect 21570 4750 30950 4760
rect 14906 3200 15086 3210
rect 14906 3120 14920 3200
rect 15070 3120 15086 3200
rect 14906 2640 15086 3120
rect 14906 2570 14920 2640
rect 15070 2570 15086 2640
rect 14906 2540 15086 2570
rect 14906 2470 14920 2540
rect 15070 2470 15086 2540
rect 14906 2459 15086 2470
rect 800 1180 1200 1190
rect 800 1110 820 1180
rect 890 1110 960 1180
rect 1030 1110 1090 1180
rect 1160 1110 1200 1180
rect 800 1080 1200 1110
rect 800 1010 820 1080
rect 890 1010 960 1080
rect 1030 1010 1090 1080
rect 1160 1010 1200 1080
rect 800 1000 1200 1010
rect 800 990 21770 1000
rect 800 920 21580 990
rect 21760 920 21770 990
rect 800 880 21770 920
rect 800 810 21580 880
rect 21760 810 21770 880
rect 800 800 21770 810
<< via3 >>
rect 27230 44950 27300 45030
rect 7920 44770 8040 44860
rect 8120 44770 8240 44860
rect 8310 44770 8430 44860
rect 27770 44880 27840 44950
rect 31460 44870 31560 44940
rect 31140 44730 31240 44800
rect 31280 44720 31380 44790
rect 31460 44760 31560 44830
rect 820 36140 910 36210
rect 960 36140 1050 36210
rect 1100 36140 1190 36210
rect 820 36020 910 36090
rect 960 36020 1050 36090
rect 1100 36020 1190 36090
rect 230 20910 300 20980
rect 350 20910 420 20980
rect 480 20910 550 20980
rect 210 20800 280 20870
rect 340 20800 410 20870
rect 470 20800 540 20870
rect 21590 4870 21750 4940
rect 30760 4870 30940 4940
rect 21590 4760 21750 4830
rect 30760 4760 30940 4830
rect 14920 3120 15070 3200
rect 14920 2570 15070 2640
rect 14920 2470 15070 2540
rect 220 1400 290 1470
rect 350 1400 420 1470
rect 480 1400 550 1470
rect 220 1290 290 1360
rect 350 1290 420 1360
rect 480 1290 550 1360
rect 820 1110 890 1180
rect 960 1110 1030 1180
rect 1090 1110 1160 1180
rect 820 1010 890 1080
rect 960 1010 1030 1080
rect 1090 1010 1160 1080
rect 21580 920 21760 990
rect 21580 810 21760 880
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 45040 27170 45152
rect 27662 45040 27722 45152
rect 27110 45030 27310 45040
rect 27110 44952 27230 45030
rect 800 44860 26647 44952
rect 27220 44950 27230 44952
rect 27300 44950 27310 45030
rect 27662 44960 27840 45040
rect 27662 44952 27850 44960
rect 27220 44940 27310 44950
rect 27760 44950 27850 44952
rect 27760 44880 27770 44950
rect 27840 44880 27850 44950
rect 28214 44938 28274 45152
rect 28766 44938 28826 45152
rect 29318 44952 29378 45152
rect 29310 44938 29378 44952
rect 27760 44870 27850 44880
rect 28210 44870 29378 44938
rect 31450 44940 31570 44950
rect 31450 44870 31460 44940
rect 31560 44870 31570 44940
rect 800 44770 7920 44860
rect 8040 44770 8120 44860
rect 8240 44770 8310 44860
rect 8430 44770 26647 44860
rect 800 44760 26647 44770
rect 28210 44760 28290 44870
rect 31450 44830 31570 44870
rect 200 20980 600 44152
rect 200 20910 230 20980
rect 300 20910 350 20980
rect 420 20910 480 20980
rect 550 20910 600 20980
rect 200 20870 600 20910
rect 200 20800 210 20870
rect 280 20800 340 20870
rect 410 20800 470 20870
rect 540 20800 600 20870
rect 200 1470 600 20800
rect 200 1400 220 1470
rect 290 1400 350 1470
rect 420 1400 480 1470
rect 550 1400 600 1470
rect 200 1360 600 1400
rect 200 1290 220 1360
rect 290 1290 350 1360
rect 420 1290 480 1360
rect 550 1290 600 1360
rect 200 1000 600 1290
rect 800 36210 1200 44760
rect 26550 44680 28290 44760
rect 31130 44800 31390 44810
rect 31130 44730 31140 44800
rect 31240 44790 31390 44800
rect 31240 44730 31280 44790
rect 31130 44720 31280 44730
rect 31380 44720 31390 44790
rect 800 36140 820 36210
rect 910 36140 960 36210
rect 1050 36140 1100 36210
rect 1190 36140 1200 36210
rect 800 36090 1200 36140
rect 800 36020 820 36090
rect 910 36020 960 36090
rect 1050 36020 1100 36090
rect 1190 36020 1200 36090
rect 800 1180 1200 36020
rect 31270 15930 31390 44720
rect 31450 44760 31460 44830
rect 31560 44760 31570 44830
rect 31450 15910 31570 44760
rect 22470 5210 22650 5520
rect 21100 5030 22650 5210
rect 800 1110 820 1180
rect 890 1110 960 1180
rect 1030 1110 1090 1180
rect 1160 1110 1200 1180
rect 800 1080 1200 1110
rect 800 1010 820 1080
rect 890 1010 960 1080
rect 1030 1010 1090 1080
rect 1160 1010 1200 1080
rect 800 1000 1200 1010
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 2990
rect 14906 2640 15086 2650
rect 14906 2570 14920 2640
rect 15070 2570 15086 2640
rect 14906 2540 15086 2570
rect 14906 2470 14920 2540
rect 15070 2470 15086 2540
rect 14906 0 15086 2470
rect 21100 1540 21280 5030
rect 18770 1360 21280 1540
rect 21570 4940 21770 4950
rect 21570 4870 21590 4940
rect 21750 4870 21770 4940
rect 21570 4830 21770 4870
rect 21570 4760 21590 4830
rect 21750 4760 21770 4830
rect 18770 0 18950 1360
rect 21570 990 21770 4760
rect 23750 4500 23930 5670
rect 21570 920 21580 990
rect 21760 920 21770 990
rect 21570 880 21770 920
rect 21570 810 21580 880
rect 21760 810 21770 880
rect 21570 800 21770 810
rect 22634 4320 23930 4500
rect 24360 4560 24540 5640
rect 30750 4940 30950 4950
rect 30750 4870 30760 4940
rect 30940 4870 30950 4940
rect 30750 4830 30950 4870
rect 30750 4760 30760 4830
rect 30940 4760 30950 4830
rect 30750 4750 30950 4760
rect 31020 4620 31200 4970
rect 24360 4380 26678 4560
rect 22634 0 22814 4320
rect 26498 0 26678 4380
rect 30362 4440 31200 4620
rect 30362 0 30542 4440
use Diff_Opamp  Diff_Opamp_0
timestamp 1757892507
transform 0 -1 31380 1 0 4920
box -3900 -190 39700 31170
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
